//this is the design file
module hello(A,B);
    input A;
    output B;
    assign B=A;
endmodule