module and_gate(A,B,C);
    input A;
    input B;
    output C;
    and(C,A,B);
endmodule