module not_gate(input A, output B);
    not(B,A);
endmodule